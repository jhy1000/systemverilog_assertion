
// Construction of sequences with temporal dealy

start ##1 transfer      // a sequence in which the boolean variable
                        // transfer holds on the clock after start.
                        
start ##2 transfer      // a sequence in which the Boolean variable 
                        // transfer holds two clocks after start.

start ##[0:2] transfer  // a sequence in which the boolean variable
                        // transfer holds between zero to two clocks
                        // after start.
