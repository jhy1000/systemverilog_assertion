

// Construction of sequences with temporal dealy

##0 a       - same as (a)
##1 a       - same as (1'b1 ##1 a)
##[0:1]     - same as a or (1'b1 ##1 a)

